 module div_by_3
(
input logic CLK,
input logic strob_RW_RD,
input logic CLR,
output logic strob_main
);






endmodule 